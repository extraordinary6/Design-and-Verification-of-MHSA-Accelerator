module lut_2D (
    input [63:0] data_in,
    input [12:0] sum,
    output [63:0] data_out
);
    
    logic [7:0] lut [1:15][1:63];
    
    initial begin
        lut[1][1] = 8'b00010000; lut[1][2] = 8'b00001000; lut[1][3] = 8'b00000101; lut[1][4] = 8'b00000100;
        lut[1][5] = 8'b00000011; lut[1][6] = 8'b00000010; lut[1][7] = 8'b00000010; lut[1][8] = 8'b00000010;
        lut[1][9] = 8'b00000001; lut[1][10] = 8'b00000001; lut[1][11] = 8'b00000001; lut[1][12] = 8'b00000001;
        lut[1][13] = 8'b00000001; lut[1][14] = 8'b00000001; lut[1][15] = 8'b00000001; lut[1][16] = 8'b00000001;
        lut[1][17] = 8'b00000000; lut[1][18] = 8'b00000000; lut[1][19] = 8'b00000000; lut[1][20] = 8'b00000000;
        lut[1][21] = 8'b00000000; lut[1][22] = 8'b00000000; lut[1][23] = 8'b00000000; lut[1][24] = 8'b00000000;
        lut[1][25] = 8'b00000000; lut[1][26] = 8'b00000000; lut[1][27] = 8'b00000000; lut[1][28] = 8'b00000000;
        lut[1][29] = 8'b00000000; lut[1][30] = 8'b00000000; lut[1][31] = 8'b00000000; lut[1][32] = 8'b00000000;
        lut[1][33] = 8'b00000000; lut[1][34] = 8'b00000000; lut[1][35] = 8'b00000000; lut[1][36] = 8'b00000000;
        lut[1][37] = 8'b00000000; lut[1][38] = 8'b00000000; lut[1][39] = 8'b00000000; lut[1][40] = 8'b00000000;
        lut[1][41] = 8'b00000000; lut[1][42] = 8'b00000000; lut[1][43] = 8'b00000000; lut[1][44] = 8'b00000000;
        lut[1][45] = 8'b00000000; lut[1][46] = 8'b00000000; lut[1][47] = 8'b00000000; lut[1][48] = 8'b00000000;
        lut[1][49] = 8'b00000000; lut[1][50] = 8'b00000000; lut[1][51] = 8'b00000000; lut[1][52] = 8'b00000000;
        lut[1][53] = 8'b00000000; lut[1][54] = 8'b00000000; lut[1][55] = 8'b00000000; lut[1][56] = 8'b00000000;
        lut[1][57] = 8'b00000000; lut[1][58] = 8'b00000000; lut[1][59] = 8'b00000000; lut[1][60] = 8'b00000000;
        lut[1][61] = 8'b00000000; lut[1][62] = 8'b00000000; lut[1][63] = 8'b00000000;
        lut[2][1] = 8'b00100000; lut[2][2] = 8'b00010000; lut[2][3] = 8'b00001010; lut[2][4] = 8'b00001000;
        lut[2][5] = 8'b00000110; lut[2][6] = 8'b00000101; lut[2][7] = 8'b00000100; lut[2][8] = 8'b00000100;
        lut[2][9] = 8'b00000011; lut[2][10] = 8'b00000011; lut[2][11] = 8'b00000010; lut[2][12] = 8'b00000010;
        lut[2][13] = 8'b00000010; lut[2][14] = 8'b00000010; lut[2][15] = 8'b00000010; lut[2][16] = 8'b00000010;
        lut[2][17] = 8'b00000001; lut[2][18] = 8'b00000001; lut[2][19] = 8'b00000001; lut[2][20] = 8'b00000001;
        lut[2][21] = 8'b00000001; lut[2][22] = 8'b00000001; lut[2][23] = 8'b00000001; lut[2][24] = 8'b00000001;
        lut[2][25] = 8'b00000001; lut[2][26] = 8'b00000001; lut[2][27] = 8'b00000001; lut[2][28] = 8'b00000001;
        lut[2][29] = 8'b00000001; lut[2][30] = 8'b00000001; lut[2][31] = 8'b00000001; lut[2][32] = 8'b00000001;
        lut[2][33] = 8'b00000000; lut[2][34] = 8'b00000000; lut[2][35] = 8'b00000000; lut[2][36] = 8'b00000000;
        lut[2][37] = 8'b00000000; lut[2][38] = 8'b00000000; lut[2][39] = 8'b00000000; lut[2][40] = 8'b00000000;
        lut[2][41] = 8'b00000000; lut[2][42] = 8'b00000000; lut[2][43] = 8'b00000000; lut[2][44] = 8'b00000000;
        lut[2][45] = 8'b00000000; lut[2][46] = 8'b00000000; lut[2][47] = 8'b00000000; lut[2][48] = 8'b00000000;
        lut[2][49] = 8'b00000000; lut[2][50] = 8'b00000000; lut[2][51] = 8'b00000000; lut[2][52] = 8'b00000000;
        lut[2][53] = 8'b00000000; lut[2][54] = 8'b00000000; lut[2][55] = 8'b00000000; lut[2][56] = 8'b00000000;
        lut[2][57] = 8'b00000000; lut[2][58] = 8'b00000000; lut[2][59] = 8'b00000000; lut[2][60] = 8'b00000000;
        lut[2][61] = 8'b00000000; lut[2][62] = 8'b00000000; lut[2][63] = 8'b00000000;
        lut[3][1] = 8'b00110000; lut[3][2] = 8'b00011000; lut[3][3] = 8'b00010000; lut[3][4] = 8'b00001100;
        lut[3][5] = 8'b00001001; lut[3][6] = 8'b00001000; lut[3][7] = 8'b00000110; lut[3][8] = 8'b00000110;
        lut[3][9] = 8'b00000101; lut[3][10] = 8'b00000100; lut[3][11] = 8'b00000100; lut[3][12] = 8'b00000100;
        lut[3][13] = 8'b00000011; lut[3][14] = 8'b00000011; lut[3][15] = 8'b00000011; lut[3][16] = 8'b00000011;
        lut[3][17] = 8'b00000010; lut[3][18] = 8'b00000010; lut[3][19] = 8'b00000010; lut[3][20] = 8'b00000010;
        lut[3][21] = 8'b00000010; lut[3][22] = 8'b00000010; lut[3][23] = 8'b00000010; lut[3][24] = 8'b00000010;
        lut[3][25] = 8'b00000001; lut[3][26] = 8'b00000001; lut[3][27] = 8'b00000001; lut[3][28] = 8'b00000001;
        lut[3][29] = 8'b00000001; lut[3][30] = 8'b00000001; lut[3][31] = 8'b00000001; lut[3][32] = 8'b00000001;
        lut[3][33] = 8'b00000001; lut[3][34] = 8'b00000001; lut[3][35] = 8'b00000001; lut[3][36] = 8'b00000001;
        lut[3][37] = 8'b00000001; lut[3][38] = 8'b00000001; lut[3][39] = 8'b00000001; lut[3][40] = 8'b00000001;
        lut[3][41] = 8'b00000001; lut[3][42] = 8'b00000001; lut[3][43] = 8'b00000001; lut[3][44] = 8'b00000001;
        lut[3][45] = 8'b00000001; lut[3][46] = 8'b00000001; lut[3][47] = 8'b00000001; lut[3][48] = 8'b00000001;
        lut[3][49] = 8'b00000000; lut[3][50] = 8'b00000000; lut[3][51] = 8'b00000000; lut[3][52] = 8'b00000000;
        lut[3][53] = 8'b00000000; lut[3][54] = 8'b00000000; lut[3][55] = 8'b00000000; lut[3][56] = 8'b00000000;
        lut[3][57] = 8'b00000000; lut[3][58] = 8'b00000000; lut[3][59] = 8'b00000000; lut[3][60] = 8'b00000000;
        lut[3][61] = 8'b00000000; lut[3][62] = 8'b00000000; lut[3][63] = 8'b00000000;
        lut[4][1] = 8'b01000000; lut[4][2] = 8'b00100000; lut[4][3] = 8'b00010101; lut[4][4] = 8'b00010000;
        lut[4][5] = 8'b00001100; lut[4][6] = 8'b00001010; lut[4][7] = 8'b00001001; lut[4][8] = 8'b00001000;
        lut[4][9] = 8'b00000111; lut[4][10] = 8'b00000110; lut[4][11] = 8'b00000101; lut[4][12] = 8'b00000101;
        lut[4][13] = 8'b00000100; lut[4][14] = 8'b00000100; lut[4][15] = 8'b00000100; lut[4][16] = 8'b00000100;
        lut[4][17] = 8'b00000011; lut[4][18] = 8'b00000011; lut[4][19] = 8'b00000011; lut[4][20] = 8'b00000011;
        lut[4][21] = 8'b00000011; lut[4][22] = 8'b00000010; lut[4][23] = 8'b00000010; lut[4][24] = 8'b00000010;
        lut[4][25] = 8'b00000010; lut[4][26] = 8'b00000010; lut[4][27] = 8'b00000010; lut[4][28] = 8'b00000010;
        lut[4][29] = 8'b00000010; lut[4][30] = 8'b00000010; lut[4][31] = 8'b00000010; lut[4][32] = 8'b00000010;
        lut[4][33] = 8'b00000001; lut[4][34] = 8'b00000001; lut[4][35] = 8'b00000001; lut[4][36] = 8'b00000001;
        lut[4][37] = 8'b00000001; lut[4][38] = 8'b00000001; lut[4][39] = 8'b00000001; lut[4][40] = 8'b00000001;
        lut[4][41] = 8'b00000001; lut[4][42] = 8'b00000001; lut[4][43] = 8'b00000001; lut[4][44] = 8'b00000001;
        lut[4][45] = 8'b00000001; lut[4][46] = 8'b00000001; lut[4][47] = 8'b00000001; lut[4][48] = 8'b00000001;
        lut[4][49] = 8'b00000001; lut[4][50] = 8'b00000001; lut[4][51] = 8'b00000001; lut[4][52] = 8'b00000001;
        lut[4][53] = 8'b00000001; lut[4][54] = 8'b00000001; lut[4][55] = 8'b00000001; lut[4][56] = 8'b00000001;
        lut[4][57] = 8'b00000001; lut[4][58] = 8'b00000001; lut[4][59] = 8'b00000001; lut[4][60] = 8'b00000001;
        lut[4][61] = 8'b00000001; lut[4][62] = 8'b00000001; lut[4][63] = 8'b00000001;
        lut[5][1] = 8'b01010000; lut[5][2] = 8'b00101000; lut[5][3] = 8'b00011010; lut[5][4] = 8'b00010100;
        lut[5][5] = 8'b00010000; lut[5][6] = 8'b00001101; lut[5][7] = 8'b00001011; lut[5][8] = 8'b00001010;
        lut[5][9] = 8'b00001000; lut[5][10] = 8'b00001000; lut[5][11] = 8'b00000111; lut[5][12] = 8'b00000110;
        lut[5][13] = 8'b00000110; lut[5][14] = 8'b00000101; lut[5][15] = 8'b00000101; lut[5][16] = 8'b00000101;
        lut[5][17] = 8'b00000100; lut[5][18] = 8'b00000100; lut[5][19] = 8'b00000100; lut[5][20] = 8'b00000100;
        lut[5][21] = 8'b00000011; lut[5][22] = 8'b00000011; lut[5][23] = 8'b00000011; lut[5][24] = 8'b00000011;
        lut[5][25] = 8'b00000011; lut[5][26] = 8'b00000011; lut[5][27] = 8'b00000010; lut[5][28] = 8'b00000010;
        lut[5][29] = 8'b00000010; lut[5][30] = 8'b00000010; lut[5][31] = 8'b00000010; lut[5][32] = 8'b00000010;
        lut[5][33] = 8'b00000010; lut[5][34] = 8'b00000010; lut[5][35] = 8'b00000010; lut[5][36] = 8'b00000010;
        lut[5][37] = 8'b00000010; lut[5][38] = 8'b00000010; lut[5][39] = 8'b00000010; lut[5][40] = 8'b00000010;
        lut[5][41] = 8'b00000001; lut[5][42] = 8'b00000001; lut[5][43] = 8'b00000001; lut[5][44] = 8'b00000001;
        lut[5][45] = 8'b00000001; lut[5][46] = 8'b00000001; lut[5][47] = 8'b00000001; lut[5][48] = 8'b00000001;
        lut[5][49] = 8'b00000001; lut[5][50] = 8'b00000001; lut[5][51] = 8'b00000001; lut[5][52] = 8'b00000001;
        lut[5][53] = 8'b00000001; lut[5][54] = 8'b00000001; lut[5][55] = 8'b00000001; lut[5][56] = 8'b00000001;
        lut[5][57] = 8'b00000001; lut[5][58] = 8'b00000001; lut[5][59] = 8'b00000001; lut[5][60] = 8'b00000001;
        lut[5][61] = 8'b00000001; lut[5][62] = 8'b00000001; lut[5][63] = 8'b00000001;
        lut[6][1] = 8'b01100000; lut[6][2] = 8'b00110000; lut[6][3] = 8'b00100000; lut[6][4] = 8'b00011000;
        lut[6][5] = 8'b00010011; lut[6][6] = 8'b00010000; lut[6][7] = 8'b00001101; lut[6][8] = 8'b00001100;
        lut[6][9] = 8'b00001010; lut[6][10] = 8'b00001001; lut[6][11] = 8'b00001000; lut[6][12] = 8'b00001000;
        lut[6][13] = 8'b00000111; lut[6][14] = 8'b00000110; lut[6][15] = 8'b00000110; lut[6][16] = 8'b00000110;
        lut[6][17] = 8'b00000101; lut[6][18] = 8'b00000101; lut[6][19] = 8'b00000101; lut[6][20] = 8'b00000100;
        lut[6][21] = 8'b00000100; lut[6][22] = 8'b00000100; lut[6][23] = 8'b00000100; lut[6][24] = 8'b00000100;
        lut[6][25] = 8'b00000011; lut[6][26] = 8'b00000011; lut[6][27] = 8'b00000011; lut[6][28] = 8'b00000011;
        lut[6][29] = 8'b00000011; lut[6][30] = 8'b00000011; lut[6][31] = 8'b00000011; lut[6][32] = 8'b00000011;
        lut[6][33] = 8'b00000010; lut[6][34] = 8'b00000010; lut[6][35] = 8'b00000010; lut[6][36] = 8'b00000010;
        lut[6][37] = 8'b00000010; lut[6][38] = 8'b00000010; lut[6][39] = 8'b00000010; lut[6][40] = 8'b00000010;
        lut[6][41] = 8'b00000010; lut[6][42] = 8'b00000010; lut[6][43] = 8'b00000010; lut[6][44] = 8'b00000010;
        lut[6][45] = 8'b00000010; lut[6][46] = 8'b00000010; lut[6][47] = 8'b00000010; lut[6][48] = 8'b00000010;
        lut[6][49] = 8'b00000001; lut[6][50] = 8'b00000001; lut[6][51] = 8'b00000001; lut[6][52] = 8'b00000001;
        lut[6][53] = 8'b00000001; lut[6][54] = 8'b00000001; lut[6][55] = 8'b00000001; lut[6][56] = 8'b00000001;
        lut[6][57] = 8'b00000001; lut[6][58] = 8'b00000001; lut[6][59] = 8'b00000001; lut[6][60] = 8'b00000001;
        lut[6][61] = 8'b00000001; lut[6][62] = 8'b00000001; lut[6][63] = 8'b00000001;
        lut[7][1] = 8'b01110000; lut[7][2] = 8'b00111000; lut[7][3] = 8'b00100101; lut[7][4] = 8'b00011100;
        lut[7][5] = 8'b00010110; lut[7][6] = 8'b00010010; lut[7][7] = 8'b00010000; lut[7][8] = 8'b00001110;
        lut[7][9] = 8'b00001100; lut[7][10] = 8'b00001011; lut[7][11] = 8'b00001010; lut[7][12] = 8'b00001001;
        lut[7][13] = 8'b00001000; lut[7][14] = 8'b00001000; lut[7][15] = 8'b00000111; lut[7][16] = 8'b00000111;
        lut[7][17] = 8'b00000110; lut[7][18] = 8'b00000110; lut[7][19] = 8'b00000101; lut[7][20] = 8'b00000101;
        lut[7][21] = 8'b00000101; lut[7][22] = 8'b00000101; lut[7][23] = 8'b00000100; lut[7][24] = 8'b00000100;
        lut[7][25] = 8'b00000100; lut[7][26] = 8'b00000100; lut[7][27] = 8'b00000100; lut[7][28] = 8'b00000100;
        lut[7][29] = 8'b00000011; lut[7][30] = 8'b00000011; lut[7][31] = 8'b00000011; lut[7][32] = 8'b00000011;
        lut[7][33] = 8'b00000011; lut[7][34] = 8'b00000011; lut[7][35] = 8'b00000011; lut[7][36] = 8'b00000011;
        lut[7][37] = 8'b00000011; lut[7][38] = 8'b00000010; lut[7][39] = 8'b00000010; lut[7][40] = 8'b00000010;
        lut[7][41] = 8'b00000010; lut[7][42] = 8'b00000010; lut[7][43] = 8'b00000010; lut[7][44] = 8'b00000010;
        lut[7][45] = 8'b00000010; lut[7][46] = 8'b00000010; lut[7][47] = 8'b00000010; lut[7][48] = 8'b00000010;
        lut[7][49] = 8'b00000010; lut[7][50] = 8'b00000010; lut[7][51] = 8'b00000010; lut[7][52] = 8'b00000010;
        lut[7][53] = 8'b00000010; lut[7][54] = 8'b00000010; lut[7][55] = 8'b00000010; lut[7][56] = 8'b00000010;
        lut[7][57] = 8'b00000001; lut[7][58] = 8'b00000001; lut[7][59] = 8'b00000001; lut[7][60] = 8'b00000001;
        lut[7][61] = 8'b00000001; lut[7][62] = 8'b00000001; lut[7][63] = 8'b00000001;
        lut[8][1] = 8'b10000000; lut[8][2] = 8'b01000000; lut[8][3] = 8'b00101010; lut[8][4] = 8'b00100000;
        lut[8][5] = 8'b00011001; lut[8][6] = 8'b00010101; lut[8][7] = 8'b00010010; lut[8][8] = 8'b00010000;
        lut[8][9] = 8'b00001110; lut[8][10] = 8'b00001100; lut[8][11] = 8'b00001011; lut[8][12] = 8'b00001010;
        lut[8][13] = 8'b00001001; lut[8][14] = 8'b00001001; lut[8][15] = 8'b00001000; lut[8][16] = 8'b00001000;
        lut[8][17] = 8'b00000111; lut[8][18] = 8'b00000111; lut[8][19] = 8'b00000110; lut[8][20] = 8'b00000110;
        lut[8][21] = 8'b00000110; lut[8][22] = 8'b00000101; lut[8][23] = 8'b00000101; lut[8][24] = 8'b00000101;
        lut[8][25] = 8'b00000101; lut[8][26] = 8'b00000100; lut[8][27] = 8'b00000100; lut[8][28] = 8'b00000100;
        lut[8][29] = 8'b00000100; lut[8][30] = 8'b00000100; lut[8][31] = 8'b00000100; lut[8][32] = 8'b00000100;
        lut[8][33] = 8'b00000011; lut[8][34] = 8'b00000011; lut[8][35] = 8'b00000011; lut[8][36] = 8'b00000011;
        lut[8][37] = 8'b00000011; lut[8][38] = 8'b00000011; lut[8][39] = 8'b00000011; lut[8][40] = 8'b00000011;
        lut[8][41] = 8'b00000011; lut[8][42] = 8'b00000011; lut[8][43] = 8'b00000010; lut[8][44] = 8'b00000010;
        lut[8][45] = 8'b00000010; lut[8][46] = 8'b00000010; lut[8][47] = 8'b00000010; lut[8][48] = 8'b00000010;
        lut[8][49] = 8'b00000010; lut[8][50] = 8'b00000010; lut[8][51] = 8'b00000010; lut[8][52] = 8'b00000010;
        lut[8][53] = 8'b00000010; lut[8][54] = 8'b00000010; lut[8][55] = 8'b00000010; lut[8][56] = 8'b00000010;
        lut[8][57] = 8'b00000010; lut[8][58] = 8'b00000010; lut[8][59] = 8'b00000010; lut[8][60] = 8'b00000010;
        lut[8][61] = 8'b00000010; lut[8][62] = 8'b00000010; lut[8][63] = 8'b00000010;
        lut[9][1] = 8'b10010000; lut[9][2] = 8'b01001000; lut[9][3] = 8'b00110000; lut[9][4] = 8'b00100100;
        lut[9][5] = 8'b00011100; lut[9][6] = 8'b00011000; lut[9][7] = 8'b00010100; lut[9][8] = 8'b00010010;
        lut[9][9] = 8'b00010000; lut[9][10] = 8'b00001110; lut[9][11] = 8'b00001101; lut[9][12] = 8'b00001100;
        lut[9][13] = 8'b00001011; lut[9][14] = 8'b00001010; lut[9][15] = 8'b00001001; lut[9][16] = 8'b00001001;
        lut[9][17] = 8'b00001000; lut[9][18] = 8'b00001000; lut[9][19] = 8'b00000111; lut[9][20] = 8'b00000111;
        lut[9][21] = 8'b00000110; lut[9][22] = 8'b00000110; lut[9][23] = 8'b00000110; lut[9][24] = 8'b00000110;
        lut[9][25] = 8'b00000101; lut[9][26] = 8'b00000101; lut[9][27] = 8'b00000101; lut[9][28] = 8'b00000101;
        lut[9][29] = 8'b00000100; lut[9][30] = 8'b00000100; lut[9][31] = 8'b00000100; lut[9][32] = 8'b00000100;
        lut[9][33] = 8'b00000100; lut[9][34] = 8'b00000100; lut[9][35] = 8'b00000100; lut[9][36] = 8'b00000100;
        lut[9][37] = 8'b00000011; lut[9][38] = 8'b00000011; lut[9][39] = 8'b00000011; lut[9][40] = 8'b00000011;
        lut[9][41] = 8'b00000011; lut[9][42] = 8'b00000011; lut[9][43] = 8'b00000011; lut[9][44] = 8'b00000011;
        lut[9][45] = 8'b00000011; lut[9][46] = 8'b00000011; lut[9][47] = 8'b00000011; lut[9][48] = 8'b00000011;
        lut[9][49] = 8'b00000010; lut[9][50] = 8'b00000010; lut[9][51] = 8'b00000010; lut[9][52] = 8'b00000010;
        lut[9][53] = 8'b00000010; lut[9][54] = 8'b00000010; lut[9][55] = 8'b00000010; lut[9][56] = 8'b00000010;
        lut[9][57] = 8'b00000010; lut[9][58] = 8'b00000010; lut[9][59] = 8'b00000010; lut[9][60] = 8'b00000010;
        lut[9][61] = 8'b00000010; lut[9][62] = 8'b00000010; lut[9][63] = 8'b00000010;
        lut[10][1] = 8'b10100000; lut[10][2] = 8'b01010000; lut[10][3] = 8'b00110101; lut[10][4] = 8'b00101000;
        lut[10][5] = 8'b00100000; lut[10][6] = 8'b00011010; lut[10][7] = 8'b00010110; lut[10][8] = 8'b00010100;
        lut[10][9] = 8'b00010001; lut[10][10] = 8'b00010000; lut[10][11] = 8'b00001110; lut[10][12] = 8'b00001101;
        lut[10][13] = 8'b00001100; lut[10][14] = 8'b00001011; lut[10][15] = 8'b00001010; lut[10][16] = 8'b00001010;
        lut[10][17] = 8'b00001001; lut[10][18] = 8'b00001000; lut[10][19] = 8'b00001000; lut[10][20] = 8'b00001000;
        lut[10][21] = 8'b00000111; lut[10][22] = 8'b00000111; lut[10][23] = 8'b00000110; lut[10][24] = 8'b00000110;
        lut[10][25] = 8'b00000110; lut[10][26] = 8'b00000110; lut[10][27] = 8'b00000101; lut[10][28] = 8'b00000101;
        lut[10][29] = 8'b00000101; lut[10][30] = 8'b00000101; lut[10][31] = 8'b00000101; lut[10][32] = 8'b00000101;
        lut[10][33] = 8'b00000100; lut[10][34] = 8'b00000100; lut[10][35] = 8'b00000100; lut[10][36] = 8'b00000100;
        lut[10][37] = 8'b00000100; lut[10][38] = 8'b00000100; lut[10][39] = 8'b00000100; lut[10][40] = 8'b00000100;
        lut[10][41] = 8'b00000011; lut[10][42] = 8'b00000011; lut[10][43] = 8'b00000011; lut[10][44] = 8'b00000011;
        lut[10][45] = 8'b00000011; lut[10][46] = 8'b00000011; lut[10][47] = 8'b00000011; lut[10][48] = 8'b00000011;
        lut[10][49] = 8'b00000011; lut[10][50] = 8'b00000011; lut[10][51] = 8'b00000011; lut[10][52] = 8'b00000011;
        lut[10][53] = 8'b00000011; lut[10][54] = 8'b00000010; lut[10][55] = 8'b00000010; lut[10][56] = 8'b00000010;
        lut[10][57] = 8'b00000010; lut[10][58] = 8'b00000010; lut[10][59] = 8'b00000010; lut[10][60] = 8'b00000010;
        lut[10][61] = 8'b00000010; lut[10][62] = 8'b00000010; lut[10][63] = 8'b00000010;
        lut[11][1] = 8'b10110000; lut[11][2] = 8'b01011000; lut[11][3] = 8'b00111010; lut[11][4] = 8'b00101100;
        lut[11][5] = 8'b00100011; lut[11][6] = 8'b00011101; lut[11][7] = 8'b00011001; lut[11][8] = 8'b00010110;
        lut[11][9] = 8'b00010011; lut[11][10] = 8'b00010001; lut[11][11] = 8'b00010000; lut[11][12] = 8'b00001110;
        lut[11][13] = 8'b00001101; lut[11][14] = 8'b00001100; lut[11][15] = 8'b00001011; lut[11][16] = 8'b00001011;
        lut[11][17] = 8'b00001010; lut[11][18] = 8'b00001001; lut[11][19] = 8'b00001001; lut[11][20] = 8'b00001000;
        lut[11][21] = 8'b00001000; lut[11][22] = 8'b00001000; lut[11][23] = 8'b00000111; lut[11][24] = 8'b00000111;
        lut[11][25] = 8'b00000111; lut[11][26] = 8'b00000110; lut[11][27] = 8'b00000110; lut[11][28] = 8'b00000110;
        lut[11][29] = 8'b00000110; lut[11][30] = 8'b00000101; lut[11][31] = 8'b00000101; lut[11][32] = 8'b00000101;
        lut[11][33] = 8'b00000101; lut[11][34] = 8'b00000101; lut[11][35] = 8'b00000101; lut[11][36] = 8'b00000100;
        lut[11][37] = 8'b00000100; lut[11][38] = 8'b00000100; lut[11][39] = 8'b00000100; lut[11][40] = 8'b00000100;
        lut[11][41] = 8'b00000100; lut[11][42] = 8'b00000100; lut[11][43] = 8'b00000100; lut[11][44] = 8'b00000100;
        lut[11][45] = 8'b00000011; lut[11][46] = 8'b00000011; lut[11][47] = 8'b00000011; lut[11][48] = 8'b00000011;
        lut[11][49] = 8'b00000011; lut[11][50] = 8'b00000011; lut[11][51] = 8'b00000011; lut[11][52] = 8'b00000011;
        lut[11][53] = 8'b00000011; lut[11][54] = 8'b00000011; lut[11][55] = 8'b00000011; lut[11][56] = 8'b00000011;
        lut[11][57] = 8'b00000011; lut[11][58] = 8'b00000011; lut[11][59] = 8'b00000010; lut[11][60] = 8'b00000010;
        lut[11][61] = 8'b00000010; lut[11][62] = 8'b00000010; lut[11][63] = 8'b00000010;
        lut[12][1] = 8'b11000000; lut[12][2] = 8'b01100000; lut[12][3] = 8'b01000000; lut[12][4] = 8'b00110000;
        lut[12][5] = 8'b00100110; lut[12][6] = 8'b00100000; lut[12][7] = 8'b00011011; lut[12][8] = 8'b00011000;
        lut[12][9] = 8'b00010101; lut[12][10] = 8'b00010011; lut[12][11] = 8'b00010001; lut[12][12] = 8'b00010000;
        lut[12][13] = 8'b00001110; lut[12][14] = 8'b00001101; lut[12][15] = 8'b00001100; lut[12][16] = 8'b00001100;
        lut[12][17] = 8'b00001011; lut[12][18] = 8'b00001010; lut[12][19] = 8'b00001010; lut[12][20] = 8'b00001001;
        lut[12][21] = 8'b00001001; lut[12][22] = 8'b00001000; lut[12][23] = 8'b00001000; lut[12][24] = 8'b00001000;
        lut[12][25] = 8'b00000111; lut[12][26] = 8'b00000111; lut[12][27] = 8'b00000111; lut[12][28] = 8'b00000110;
        lut[12][29] = 8'b00000110; lut[12][30] = 8'b00000110; lut[12][31] = 8'b00000110; lut[12][32] = 8'b00000110;
        lut[12][33] = 8'b00000101; lut[12][34] = 8'b00000101; lut[12][35] = 8'b00000101; lut[12][36] = 8'b00000101;
        lut[12][37] = 8'b00000101; lut[12][38] = 8'b00000101; lut[12][39] = 8'b00000100; lut[12][40] = 8'b00000100;
        lut[12][41] = 8'b00000100; lut[12][42] = 8'b00000100; lut[12][43] = 8'b00000100; lut[12][44] = 8'b00000100;
        lut[12][45] = 8'b00000100; lut[12][46] = 8'b00000100; lut[12][47] = 8'b00000100; lut[12][48] = 8'b00000100;
        lut[12][49] = 8'b00000011; lut[12][50] = 8'b00000011; lut[12][51] = 8'b00000011; lut[12][52] = 8'b00000011;
        lut[12][53] = 8'b00000011; lut[12][54] = 8'b00000011; lut[12][55] = 8'b00000011; lut[12][56] = 8'b00000011;
        lut[12][57] = 8'b00000011; lut[12][58] = 8'b00000011; lut[12][59] = 8'b00000011; lut[12][60] = 8'b00000011;
        lut[12][61] = 8'b00000011; lut[12][62] = 8'b00000011; lut[12][63] = 8'b00000011;
        lut[13][1] = 8'b11010000; lut[13][2] = 8'b01101000; lut[13][3] = 8'b01000101; lut[13][4] = 8'b00110100;
        lut[13][5] = 8'b00101001; lut[13][6] = 8'b00100010; lut[13][7] = 8'b00011101; lut[13][8] = 8'b00011010;
        lut[13][9] = 8'b00010111; lut[13][10] = 8'b00010100; lut[13][11] = 8'b00010010; lut[13][12] = 8'b00010001;
        lut[13][13] = 8'b00010000; lut[13][14] = 8'b00001110; lut[13][15] = 8'b00001101; lut[13][16] = 8'b00001101;
        lut[13][17] = 8'b00001100; lut[13][18] = 8'b00001011; lut[13][19] = 8'b00001010; lut[13][20] = 8'b00001010;
        lut[13][21] = 8'b00001001; lut[13][22] = 8'b00001001; lut[13][23] = 8'b00001001; lut[13][24] = 8'b00001000;
        lut[13][25] = 8'b00001000; lut[13][26] = 8'b00001000; lut[13][27] = 8'b00000111; lut[13][28] = 8'b00000111;
        lut[13][29] = 8'b00000111; lut[13][30] = 8'b00000110; lut[13][31] = 8'b00000110; lut[13][32] = 8'b00000110;
        lut[13][33] = 8'b00000110; lut[13][34] = 8'b00000110; lut[13][35] = 8'b00000101; lut[13][36] = 8'b00000101;
        lut[13][37] = 8'b00000101; lut[13][38] = 8'b00000101; lut[13][39] = 8'b00000101; lut[13][40] = 8'b00000101;
        lut[13][41] = 8'b00000101; lut[13][42] = 8'b00000100; lut[13][43] = 8'b00000100; lut[13][44] = 8'b00000100;
        lut[13][45] = 8'b00000100; lut[13][46] = 8'b00000100; lut[13][47] = 8'b00000100; lut[13][48] = 8'b00000100;
        lut[13][49] = 8'b00000100; lut[13][50] = 8'b00000100; lut[13][51] = 8'b00000100; lut[13][52] = 8'b00000100;
        lut[13][53] = 8'b00000011; lut[13][54] = 8'b00000011; lut[13][55] = 8'b00000011; lut[13][56] = 8'b00000011;
        lut[13][57] = 8'b00000011; lut[13][58] = 8'b00000011; lut[13][59] = 8'b00000011; lut[13][60] = 8'b00000011;
        lut[13][61] = 8'b00000011; lut[13][62] = 8'b00000011; lut[13][63] = 8'b00000011;
        lut[14][1] = 8'b11100000; lut[14][2] = 8'b01110000; lut[14][3] = 8'b01001010; lut[14][4] = 8'b00111000;
        lut[14][5] = 8'b00101100; lut[14][6] = 8'b00100101; lut[14][7] = 8'b00100000; lut[14][8] = 8'b00011100;
        lut[14][9] = 8'b00011000; lut[14][10] = 8'b00010110; lut[14][11] = 8'b00010100; lut[14][12] = 8'b00010010;
        lut[14][13] = 8'b00010001; lut[14][14] = 8'b00010000; lut[14][15] = 8'b00001110; lut[14][16] = 8'b00001110;
        lut[14][17] = 8'b00001101; lut[14][18] = 8'b00001100; lut[14][19] = 8'b00001011; lut[14][20] = 8'b00001011;
        lut[14][21] = 8'b00001010; lut[14][22] = 8'b00001010; lut[14][23] = 8'b00001001; lut[14][24] = 8'b00001001;
        lut[14][25] = 8'b00001000; lut[14][26] = 8'b00001000; lut[14][27] = 8'b00001000; lut[14][28] = 8'b00001000;
        lut[14][29] = 8'b00000111; lut[14][30] = 8'b00000111; lut[14][31] = 8'b00000111; lut[14][32] = 8'b00000111;
        lut[14][33] = 8'b00000110; lut[14][34] = 8'b00000110; lut[14][35] = 8'b00000110; lut[14][36] = 8'b00000110;
        lut[14][37] = 8'b00000110; lut[14][38] = 8'b00000101; lut[14][39] = 8'b00000101; lut[14][40] = 8'b00000101;
        lut[14][41] = 8'b00000101; lut[14][42] = 8'b00000101; lut[14][43] = 8'b00000101; lut[14][44] = 8'b00000101;
        lut[14][45] = 8'b00000100; lut[14][46] = 8'b00000100; lut[14][47] = 8'b00000100; lut[14][48] = 8'b00000100;
        lut[14][49] = 8'b00000100; lut[14][50] = 8'b00000100; lut[14][51] = 8'b00000100; lut[14][52] = 8'b00000100;
        lut[14][53] = 8'b00000100; lut[14][54] = 8'b00000100; lut[14][55] = 8'b00000100; lut[14][56] = 8'b00000100;
        lut[14][57] = 8'b00000011; lut[14][58] = 8'b00000011; lut[14][59] = 8'b00000011; lut[14][60] = 8'b00000011;
        lut[14][61] = 8'b00000011; lut[14][62] = 8'b00000011; lut[14][63] = 8'b00000011;
        lut[15][1] = 8'b11110000; lut[15][2] = 8'b01111000; lut[15][3] = 8'b01010000; lut[15][4] = 8'b00111100;
        lut[15][5] = 8'b00110000; lut[15][6] = 8'b00101000; lut[15][7] = 8'b00100010; lut[15][8] = 8'b00011110;
        lut[15][9] = 8'b00011010; lut[15][10] = 8'b00011000; lut[15][11] = 8'b00010101; lut[15][12] = 8'b00010100;
        lut[15][13] = 8'b00010010; lut[15][14] = 8'b00010001; lut[15][15] = 8'b00010000; lut[15][16] = 8'b00001111;
        lut[15][17] = 8'b00001110; lut[15][18] = 8'b00001101; lut[15][19] = 8'b00001100; lut[15][20] = 8'b00001100;
        lut[15][21] = 8'b00001011; lut[15][22] = 8'b00001010; lut[15][23] = 8'b00001010; lut[15][24] = 8'b00001010;
        lut[15][25] = 8'b00001001; lut[15][26] = 8'b00001001; lut[15][27] = 8'b00001000; lut[15][28] = 8'b00001000;
        lut[15][29] = 8'b00001000; lut[15][30] = 8'b00001000; lut[15][31] = 8'b00000111; lut[15][32] = 8'b00000111;
        lut[15][33] = 8'b00000111; lut[15][34] = 8'b00000111; lut[15][35] = 8'b00000110; lut[15][36] = 8'b00000110;
        lut[15][37] = 8'b00000110; lut[15][38] = 8'b00000110; lut[15][39] = 8'b00000110; lut[15][40] = 8'b00000110;
        lut[15][41] = 8'b00000101; lut[15][42] = 8'b00000101; lut[15][43] = 8'b00000101; lut[15][44] = 8'b00000101;
        lut[15][45] = 8'b00000101; lut[15][46] = 8'b00000101; lut[15][47] = 8'b00000101; lut[15][48] = 8'b00000101;
        lut[15][49] = 8'b00000100; lut[15][50] = 8'b00000100; lut[15][51] = 8'b00000100; lut[15][52] = 8'b00000100;
        lut[15][53] = 8'b00000100; lut[15][54] = 8'b00000100; lut[15][55] = 8'b00000100; lut[15][56] = 8'b00000100;
        lut[15][57] = 8'b00000100; lut[15][58] = 8'b00000100; lut[15][59] = 8'b00000100; lut[15][60] = 8'b00000100;
        lut[15][61] = 8'b00000011; lut[15][62] = 8'b00000011; lut[15][63] = 8'b00000011;
    end

    logic [5:0] sum_p;
        
    assign sum_p = sum[12:7];

    assign data_out[7:0] = (data_in[7:0] != 0 && sum_p != 0) ? lut[data_in[7:4]][sum_p] : 0;
    assign data_out[15:8] = (data_in[15:8] != 0 && sum_p != 0) ? lut[data_in[15:12]][sum_p] : 0;
    assign data_out[23:16] = (data_in[23:16] != 0 && sum_p != 0) ? lut[data_in[23:20]][sum_p] : 0;
    assign data_out[31:24] = (data_in[31:24] != 0 && sum_p != 0) ? lut[data_in[31:28]][sum_p] : 0;
    assign data_out[39:32] = (data_in[39:32] != 0 && sum_p != 0) ? lut[data_in[39:36]][sum_p] : 0;
    assign data_out[47:40] = (data_in[47:40] != 0 && sum_p != 0) ? lut[data_in[47:44]][sum_p] : 0;
    assign data_out[55:48] = (data_in[55:48] != 0 && sum_p != 0) ? lut[data_in[55:52]][sum_p] : 0;
    assign data_out[63:56] = (data_in[63:56] != 0 && sum_p != 0) ? lut[data_in[63:60]][sum_p] : 0;

endmodule