module lut_1D (
    input [63:0] data_in,
    output [63:0] data_out
);
    
    logic [7:0] lut [0:255];
    
    // data_in / (64 + 32)
    initial begin
        lut[0] = 8'b00010001; lut[1] = 8'b00010010; lut[2] = 8'b00010010; lut[3] = 8'b00010010;
        lut[4] = 8'b00010010; lut[5] = 8'b00010010; lut[6] = 8'b00010011; lut[7] = 8'b00010011;
        lut[8] = 8'b00010011; lut[9] = 8'b00010011; lut[10] = 8'b00010011; lut[11] = 8'b00010100;
        lut[12] = 8'b00010100; lut[13] = 8'b00010100; lut[14] = 8'b00010100; lut[15] = 8'b00010100;
        lut[16] = 8'b00010101; lut[17] = 8'b00010101; lut[18] = 8'b00010101; lut[19] = 8'b00010101;
        lut[20] = 8'b00010110; lut[21] = 8'b00010110; lut[22] = 8'b00010110; lut[23] = 8'b00010110;
        lut[24] = 8'b00010110; lut[25] = 8'b00010111; lut[26] = 8'b00010111; lut[27] = 8'b00010111;
        lut[28] = 8'b00010111; lut[29] = 8'b00011000; lut[30] = 8'b00011000; lut[31] = 8'b00011000;
        lut[32] = 8'b00011000; lut[33] = 8'b00011001; lut[34] = 8'b00011001; lut[35] = 8'b00011001;
        lut[36] = 8'b00011010; lut[37] = 8'b00011010; lut[38] = 8'b00011010; lut[39] = 8'b00011010;
        lut[40] = 8'b00011011; lut[41] = 8'b00011011; lut[42] = 8'b00011011; lut[43] = 8'b00011100;
        lut[44] = 8'b00011100; lut[45] = 8'b00011100; lut[46] = 8'b00011100; lut[47] = 8'b00011101;
        lut[48] = 8'b00011101; lut[49] = 8'b00011101; lut[50] = 8'b00011110; lut[51] = 8'b00011110;
        lut[52] = 8'b00011110; lut[53] = 8'b00011111; lut[54] = 8'b00011111; lut[55] = 8'b00011111;
        lut[56] = 8'b00100000; lut[57] = 8'b00100000; lut[58] = 8'b00100000; lut[59] = 8'b00100001;
        lut[60] = 8'b00100001; lut[61] = 8'b00100001; lut[62] = 8'b00100010; lut[63] = 8'b00100010;
        lut[64] = 8'b00100010; lut[65] = 8'b00100011; lut[66] = 8'b00100011; lut[67] = 8'b00100011;
        lut[68] = 8'b00100100; lut[69] = 8'b00100100; lut[70] = 8'b00100101; lut[71] = 8'b00100101;
        lut[72] = 8'b00100101; lut[73] = 8'b00100110; lut[74] = 8'b00100110; lut[75] = 8'b00100111;
        lut[76] = 8'b00100111; lut[77] = 8'b00100111; lut[78] = 8'b00101000; lut[79] = 8'b00101000;
        lut[80] = 8'b00101001; lut[81] = 8'b00101001; lut[82] = 8'b00101010; lut[83] = 8'b00101010;
        lut[84] = 8'b00101010; lut[85] = 8'b00101011; lut[86] = 8'b00101011; lut[87] = 8'b00101100;
        lut[88] = 8'b00101100; lut[89] = 8'b00101101; lut[90] = 8'b00101101; lut[91] = 8'b00101110;
        lut[92] = 8'b00101110; lut[93] = 8'b00101111; lut[94] = 8'b00101111; lut[95] = 8'b00110000;
        lut[96] = 8'b00110000; lut[97] = 8'b00110001; lut[98] = 8'b00110001; lut[99] = 8'b00110010;
        lut[100] = 8'b00110010; lut[101] = 8'b00110011; lut[102] = 8'b00110011; lut[103] = 8'b00110100;
        lut[104] = 8'b00110100; lut[105] = 8'b00110101; lut[106] = 8'b00110110; lut[107] = 8'b00110110;
        lut[108] = 8'b00110111; lut[109] = 8'b00110111; lut[110] = 8'b00111000; lut[111] = 8'b00111000;
        lut[112] = 8'b00111001; lut[113] = 8'b00111010; lut[114] = 8'b00111010; lut[115] = 8'b00111011;
        lut[116] = 8'b00111011; lut[117] = 8'b00111100; lut[118] = 8'b00111101; lut[119] = 8'b00111101;
        lut[120] = 8'b00111110; lut[121] = 8'b00111111; lut[122] = 8'b00111111; lut[123] = 8'b01000000;
        lut[124] = 8'b01000001; lut[125] = 8'b01000001; lut[126] = 8'b01000010; lut[127] = 8'b01000011;
        lut[128] = 8'b01000011; lut[129] = 8'b01000100; lut[130] = 8'b01000101; lut[131] = 8'b01000110;
        lut[132] = 8'b01000110; lut[133] = 8'b01000111; lut[134] = 8'b01001000; lut[135] = 8'b01001001;
        lut[136] = 8'b01001001; lut[137] = 8'b01001010; lut[138] = 8'b01001011; lut[139] = 8'b01001100;
        lut[140] = 8'b01001100; lut[141] = 8'b01001101; lut[142] = 8'b01001110; lut[143] = 8'b01001111;
        lut[144] = 8'b01010000; lut[145] = 8'b01010001; lut[146] = 8'b01010001; lut[147] = 8'b01010010;
        lut[148] = 8'b01010011; lut[149] = 8'b01010100; lut[150] = 8'b01010101; lut[151] = 8'b01010110;
        lut[152] = 8'b01010111; lut[153] = 8'b01011000; lut[154] = 8'b01011001; lut[155] = 8'b01011001;
        lut[156] = 8'b01011010; lut[157] = 8'b01011011; lut[158] = 8'b01011100; lut[159] = 8'b01011101;
        lut[160] = 8'b01011110; lut[161] = 8'b01011111; lut[162] = 8'b01100000; lut[163] = 8'b01100001;
        lut[164] = 8'b01100010; lut[165] = 8'b01100011; lut[166] = 8'b01100100; lut[167] = 8'b01100101;
        lut[168] = 8'b01100111; lut[169] = 8'b01101000; lut[170] = 8'b01101001; lut[171] = 8'b01101010;
        lut[172] = 8'b01101011; lut[173] = 8'b01101100; lut[174] = 8'b01101101; lut[175] = 8'b01101110;
        lut[176] = 8'b01101111; lut[177] = 8'b01110001; lut[178] = 8'b01110010; lut[179] = 8'b01110011;
        lut[180] = 8'b01110100; lut[181] = 8'b01110101; lut[182] = 8'b01110111; lut[183] = 8'b01111000;
        lut[184] = 8'b01111001; lut[185] = 8'b01111010; lut[186] = 8'b01111100; lut[187] = 8'b01111101;
        lut[188] = 8'b01111110; lut[189] = 8'b10000000; lut[190] = 8'b10000001; lut[191] = 8'b10000010;
        lut[192] = 8'b10000100; lut[193] = 8'b10000101; lut[194] = 8'b10000111; lut[195] = 8'b10001000;
        lut[196] = 8'b10001001; lut[197] = 8'b10001011; lut[198] = 8'b10001100; lut[199] = 8'b10001110;
        lut[200] = 8'b10001111; lut[201] = 8'b10010001; lut[202] = 8'b10010010; lut[203] = 8'b10010100;
        lut[204] = 8'b10010101; lut[205] = 8'b10010111; lut[206] = 8'b10011001; lut[207] = 8'b10011010;
        lut[208] = 8'b10011100; lut[209] = 8'b10011101; lut[210] = 8'b10011111; lut[211] = 8'b10100001;
        lut[212] = 8'b10100010; lut[213] = 8'b10100100; lut[214] = 8'b10100110; lut[215] = 8'b10101000;
        lut[216] = 8'b10101001; lut[217] = 8'b10101011; lut[218] = 8'b10101101; lut[219] = 8'b10101111;
        lut[220] = 8'b10110001; lut[221] = 8'b10110010; lut[222] = 8'b10110100; lut[223] = 8'b10110110;
        lut[224] = 8'b10111000; lut[225] = 8'b10111010; lut[226] = 8'b10111100; lut[227] = 8'b10111110;
        lut[228] = 8'b11000000; lut[229] = 8'b11000010; lut[230] = 8'b11000100; lut[231] = 8'b11000110;
        lut[232] = 8'b11001000; lut[233] = 8'b11001010; lut[234] = 8'b11001100; lut[235] = 8'b11001111;
        lut[236] = 8'b11010001; lut[237] = 8'b11010011; lut[238] = 8'b11010101; lut[239] = 8'b11010111;
        lut[240] = 8'b11011010; lut[241] = 8'b11011100; lut[242] = 8'b11011110; lut[243] = 8'b11100001;
        lut[244] = 8'b11100011; lut[245] = 8'b11100101; lut[246] = 8'b11101000; lut[247] = 8'b11101010;
        lut[248] = 8'b11101101; lut[249] = 8'b11101111; lut[250] = 8'b11110010; lut[251] = 8'b11110100;
        lut[252] = 8'b11110111; lut[253] = 8'b11111001; lut[254] = 8'b11111100; lut[255] = 8'b11111111;
    end
    
    assign data_out[7:0] = lut[data_in[7:0]];
    assign data_out[15:8] = lut[data_in[15:8]];
    assign data_out[23:16] = lut[data_in[23:16]];
    assign data_out[31:24] = lut[data_in[31:24]];
    assign data_out[39:32] = lut[data_in[39:32]];
    assign data_out[47:40] = lut[data_in[47:40]];
    assign data_out[55:48] = lut[data_in[55:48]];
    assign data_out[63:56] = lut[data_in[63:56]];

endmodule