//===================================================================== 
// Description: 
// soc icb to usram bus interface, 32bit to 64bit
// Designer : wangziyao1@sjtu.edu.cn
// Revision History: 
// V0 date:Initial version @ 2024/4/21
// ==================================================================== 

// ��SOC���Բ���ͳһ��ַ�ռ䣬��ÿ��bar�ĵ�ַ�������ص�